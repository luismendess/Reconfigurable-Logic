library ieee;
use ieee.numeric_std.all;

package my_types_pkg is
    type unsigned_array is array (natural range <>) of unsigned;
end package my_types_pkg;